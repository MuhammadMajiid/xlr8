library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity char_rom is
    port (
        ascii_char : in std_logic_vector (6 downto 0);
        gdram_char : out std_logic_vector (63 downto 0)
    );
end entity;

architecture rtl of char_rom is
type GDRAM is array (0 to 127) of std_logic_vector (63 downto 0);
constant ram : GDRAM := (
    0 => x"0000000000000000",
    1 => x"0000000000000000",
    2 => x"0000000000000000",
    3 => x"0000000000000000",
    4 => x"0000000000000000",
    5 => x"0000000000000000",
    6 => x"0000000000000000",
    7 => x"0000000000000000",
    8 => x"0000000000000000",
    9 => x"0000000000000000",
    10 => x"0000000000000000",
    11 => x"0000000000000000",
    12 => x"0000000000000000",
    13 => x"0000000000000000",
    14 => x"0000000000000000",
    15 => x"0000000000000000",
    16 => x"0000000000000000",
    17 => x"0000000000000000",
    18 => x"0000000000000000",
    19 => x"0000000000000000",
    20 => x"0000000000000000",
    21 => x"0000000000000000",
    22 => x"0000000000000000",
    23 => x"0000000000000000",
    24 => x"0000000000000000",
    25 => x"0000000000000000",
    26 => x"0000000000000000",
    27 => x"0000000000000000",
    28 => x"0000000000000000",
    29 => x"0000000000000000",
    30 => x"0000000000000000",
    31 => x"0000000000000000",
    32 => x"0000000000000000",
    33 => x"0000005f00000000",--    !
    34 => x"0000030003000000",--    "
    35 => x"643c26643c262400",--    #
    36 => x"2649497f49493200",--    $
    37 => x"4225120824522100",--    %
    38 => x"20504e5522582800",--    &
    39 => x"0000000300000000",--    '
    40 => x"00001c2241000000",--    (
    41 => x"00000041221c0000",--    )
    42 => x"0015150e0e151500",--    *
    43 => x"0008083e08080000",--    +
    44 => x"0000005030000000",--    ,
    45 => x"0008080808080000",--    -
    46 => x"0000004000000000",--    .
    47 => x"4020100804020100",--    /
    48 => x"003e4141413e0000",--    0
    49 => x"0000417f40000000",--    1
    50 => x"00426151496e0000",--    2
    51 => x"0022414949360000",--    3
    52 => x"001814127f100000",--    4
    53 => x"0027494949710000",--    5
    54 => x"003c4a4948700000",--    6
    55 => x"004321110d030000",--    7
    56 => x"0036494949360000",--    8
    57 => x"00060949291e0000",--    9
    58 => x"0000001200000000",--    :
    59 => x"0000005230000000",--    ;
    60 => x"0000081414220000",--    <
    61 => x"0014141414141400",--    =
    62 => x"0000221414080000",--    >
    63 => x"0002015905020000",--    ?
    64 => x"3e415d554d512e00",--    @
    65 => x"407c4a094a7c4000",--    A
    66 => x"417f494949493600",--    B
    67 => x"1c22414141412200",--    C
    68 => x"417f414141221c00",--    D
    69 => x"417f49495d416300",--    E
    70 => x"417f49091d010300",--    F
    71 => x"1c224149493a0800",--    G
    72 => x"417f0808087f4100",--    H
    73 => x"0041417f41410000",--    I
    74 => x"304041413f010100",--    J
    75 => x"417f080c12614100",--    K
    76 => x"417f414040406000",--    L
    77 => x"417f420c427f4100",--    M
    78 => x"417f420c117f0100",--    N
    79 => x"1c22414141221c00",--    O
    80 => x"417f490909090600",--    P
    81 => x"0c12212161524c00",--    Q
    82 => x"417f090919694600",--    R
    83 => x"6649494949493300",--    S
    84 => x"0301417f41010300",--    T
    85 => x"013f4140413f0100",--    U
    86 => x"010f3140310f0100",--    V
    87 => x"011f6114611f0100",--    W
    88 => x"4141360836414100",--    X
    89 => x"0103447844030100",--    Y
    90 => x"4361514945436100",--    Z
    91 => x"00007f4141000000",--    [
    92 => x"0102040810204000",--    \
    93 => x"000041417f000000",--    ]
    94 => x"0004020101020400",--    ^
    95 => x"0040404040404000",--    _
    96 => x"0001020000000000",--    `
    97 => x"00344a4a4a3c4000",--    a
    98 => x"00413f4848483000",--    b
    99 => x"003c424242240000",--    c
    100 => x"00304848493f4000",--    d
    101 => x"003c4a4a4a2c0000",--    e
    102 => x"0000487e49090000",--    f
    103 => x"00264949493f0100",--    g
    104 => x"417f480444784000",--    h
    105 => x"0000447d40000000",--    i
    106 => x"000040443d000000",--    j
    107 => x"417f101824424200",--    k
    108 => x"0040417f40400000",--    l
    109 => x"427e027c027e4000",--    m
    110 => x"427e4402427c4000",--    n
    111 => x"003c4242423c0000",--    o
    112 => x"00417f4909090600",--    p
    113 => x"00060909497f4100",--    q
    114 => x"00427e4402020400",--    r
    115 => x"00644a4a4a360000",--    s
    116 => x"00043f4444200000",--    t
    117 => x"00023e4040227e40",--    u
    118 => x"020e3240320e0200",--    v
    119 => x"021e6218621e0200",--    w
    120 => x"4262140814624200",--    x
    121 => x"0143453805030100",--    y
    122 => x"004662524a466200",--    z
    123 => x"0000083641000000",--    {
    124 => x"0000007f00000000",--    |
    125 => x"0000004136080000",--    }
    126 => x"0018080810101800",--    ~
    127 => x"aa55aa55aa55aa55"--    DEL
); 
begin
    gdram_char <= ram(to_integer(unsigned(ascii_char)));
end architecture;